LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;
-----------------------------------------------------
ENTITY uProgramMemory IS
PORT(	
		uaddr	:	IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
		U_I	: 	OUT 	STD_LOGIC_VECTOR(28 DOWNTO 0));
END ENTITY uProgramMemory;
-----------------------------------------------------
ARCHITECTURE behavioral OF uProgramMemory IS
BEGIN
	
	MU_I: PROCESS(uaddr) 
	BEGIN
		CASE uaddr IS
	
			-- FETCH 							    
			WHEN "00000000" => U_I <= "00000000000100000000010110100"; 
			WHEN "00000001" => U_I <= "00000010000000000000010000000"; 
			WHEN "00000010" => U_I <= "00110001000000010000010000000"; 
			WHEN "00000011" => U_I <= "00000100000000100000001000000"; 
																					
			-- INT
			WHEN "00000100" => U_I <= "00000000000000000000110000000"; 
 

			--00001	 MOV ACC,A 
			WHEN "00001000" => U_I <= "00000001111011000101001000000";
       
			--00010  MOV A,ACC
			WHEN "00010000" => U_I <= "00000001011111000101111000000";
			
			
			--00011	 MOV ACC,CTE
			WHEN "00011000" => U_I <= "00000010000000000000010000000";
			
			
			--00100  MOV ACC,[DPTR]
			WHEN "00100000" => U_I <= "00000010000010000000010000000";
			

			--00101  MOV DPTR,ACC
			WHEN "00101000" => U_I <= "00000001010111000100000000000";
		
			
			-- 00110 MOV [DPTR],ACC	
			WHEN "00110000" => U_I <= "00000010000010000011101000000";
	  

			-- 00111 INV ACC
			WHEN "00111000" => U_I <= "00001010000000000100000000000";
		
			 -- 01000 AND ACC,A	 
			WHEN "01000000" => U_I <= "00000001010100000100000000000";

			
			-- 01001 ADD ACC,A
			WHEN "01001000" => U_I <= "00101001111011000100000000000";
	
			
			-- 01010 JMP DIR
			WHEN "01010000" => U_I <= "00000010000000000011111001000";
			WHEN "01010001" => U_I <= "00110001000000010011111000000";
			WHEN "01010010" => U_I <= "00000010001000000010000000000";
	
			
			-- 01011 JZ DIR
			WHEN "01011000" => U_I <= "00000000000000000001111001000";
			WHEN "01011001" => U_I <= "00000001010000000000000000000";
			WHEN "01011010" => U_I <= "00000010000010000011111000000";
			WHEN "01011011" => U_I <= "00000100001000110010000000000";
		
			
			-- 01100 JN DIR
			WHEN "01100000" => U_I <= "00000000000000000001111011000";
			WHEN "01100001" => U_I <= "00000100000000100000001000000";
			WHEN "01100010" => U_I <= "00000010000001000011111000000";
			WHEN "01100011" => U_I <= "00000100001000110010000000000";
			
			
			-- 01101 JC DIR
			WHEN "01101000" => U_I <= "00000000000000000000010100010";
			WHEN "01101001" => U_I <= "00110001000000000001000000000";
			WHEN "01101010" => U_I <= "00000010000000000000010000000";
			WHEN "01101011" => U_I <= "00000000000000110000010000000";
			WHEN "01101100" => U_I <= "00000001000000010001001000000";
			
			
			-- 01110  CALL DIR       
			WHEN "01110000" => U_I <= "00000010000001000011111000000";
			WHEN "01110001" => U_I <= "00000001001100010011111000000";
			WHEN "01110010" => U_I <= "00000001001001000011111000000";
			WHEN "01110011" => U_I <= "00000010000001000011111000000";
			WHEN "01110100" => U_I <= "00000000000001111011111000000";
			WHEN "01110101" => U_I <= "00000001000010000011111000000";
		
			
			
			-- 01111  RET
			WHEN "01111000" => U_I <= "00000001110111000001111000000";
			WHEN "01111001" => U_I <= "00000001111010000001111000000";
			WHEN "01111010" => U_I <= "00000001010110000001111000000";
			WHEN "01111011" => U_I <= "00000010000010000011111000000";
			WHEN "01111100" => U_I <= "00000001001000110011111000000";
			WHEN "01111101" => U_I <= "00000001111101000000000000000";
			
			
		
	    
	

			WHEN others => U_I <= (others => 'X');
		END CASE;
	END PROCESS;
END ARCHITECTURE Behavioral;




